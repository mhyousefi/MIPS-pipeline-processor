class generator; 

